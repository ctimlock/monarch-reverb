* C:\Users\Charlie\Projects\amp-work\Benson Monarch\LTSpice\HammondTransformer.asc
l�p1 p1 n006 5 rser=12.46 
r:u1:swa12 p2 n005 0.001 
r:u1:swa13 p2 p1 1000000000000 
r:u1:swa23 n005 p1 1000000000000 
r:u1:swb12 n006 n005 0.001 
r:u1:swb13 n006 - 1000000000000 
r:u1:swb23 n005 - 1000000000000 
l�hv1 n002 n001 22.1375868055556 rser=132.211538461539 
l�hv2 n003 n002 0.875013888888889 rser=0.961538461538407 
l�hv3 n004 n003 31.81503125 rser=133.173076923077 
l�rf1 n008 n007 0.00268154201388888 rser=0.0697499999999991 
l�rf2 n009 n008 0.00268154201388888 rser=0.0697499999999991 
l�ht1 n011 n010 0.004343878125 rser=0.0645 
l�ht2 n012 n011 0.004343878125 rser=0.0645 
l�p2 p2 - 5 rser=12.46 
k1_A0 p1 p2 0.995
k1_A1 p1 hv1 0.995
k1_A2 p1 hv2 0.995
k1_A3 p1 hv3 0.995
k1_A4 p1 rf1 0.995
k1_A5 p1 rf2 0.995
k1_A6 p1 ht1 0.995
k1_A7 p1 ht2 0.995
k1_A8 p2 hv1 0.995
k1_A9 p2 hv2 0.995
k1_A10 p2 hv3 0.995
k1_A11 p2 rf1 0.995
k1_A12 p2 rf2 0.995
k1_A13 p2 ht1 0.995
k1_A14 p2 ht2 0.995
k1_A15 hv1 hv2 0.995
k1_A16 hv1 hv3 0.995
k1_A17 hv1 rf1 0.995
k1_A18 hv1 rf2 0.995
k1_A19 hv1 ht1 0.995
k1_A20 hv1 ht2 0.995
k1_A21 hv2 hv3 0.995
k1_A22 hv2 rf1 0.995
k1_A23 hv2 rf2 0.995
k1_A24 hv2 ht1 0.995
k1_A25 hv2 ht2 0.995
k1_A26 hv3 rf1 0.995
k1_A27 hv3 rf2 0.995
k1_A28 hv3 ht1 0.995
k1_A29 hv3 ht2 0.995
k1_A30 rf1 rf2 0.995
k1_A31 rf1 ht1 0.995
k1_A32 rf1 ht2 0.995
k1_A33 rf2 ht1 0.995
k1_A34 rf2 ht2 0.995
k1_A35 ht1 ht2 0.995
.tran 0 1 0
.end
